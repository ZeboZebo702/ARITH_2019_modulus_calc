module x_500_mod_4051(
    input [500:1] X,
    output [12:1] R
    );

wire [29:1] R_temp_1;
wire [18:1] R_temp_2;
wire [13:1] R_temp_3;
wire [13:1] R_temp_4;
reg [12:1]  R_temp;

assign R_temp_1 = X [ 12 : 1 ]  + X [ 24 : 13 ] * 6'b101101 + X [ 36 : 25 ] * 11'b11111101001 + 
						X [ 48 : 37 ] * 11'b11111010011 + X [ 60 : 49 ] * 10'b1111110101 + 
						X [ 72 : 61 ] * 11'b10000000000 + X [ 84 : 73 ] * 11'b10111101111 + 
						X [ 96 : 85 ] * 12'b110111010011 + X [ 108 : 97 ] * 11'b10011110010 + 
						X [ 120 : 109 ] * 9'b100000000 + X [ 132 : 121 ] * 12'b110101011010 + 
						X [ 144 : 133 ] * 12'b111101010011 + X [ 156 : 145 ] * 12'b100100100110 + 
						{X [ 168 : 157 ], 6'b000000} + X [ 180 : 169 ] * 12'b101101000000 + 
						X [ 192 : 181 ] * 12'b111110110011 + X [ 204 : 193 ] * 12'b101000110011 + 
						{X [ 216 : 205 ], 4'b0000} + X [ 228 : 217 ] * 10'b1011010000 + 
						X [ 240 : 229 ] * 12'b111111001011 + X [ 252 : 241 ] * 12'b111001101011 + 
						{X [ 264 : 253 ], 2'b00} + X [ 276 : 265 ] * 8'b10110100 + 
						X [ 288 : 277 ] * 12'b111111010001 + X [ 300 : 289 ] * 12'b111101111001 + 
						X [ 312 : 301 ]  + X [ 324 : 313 ] * 6'b101101 + X [ 336 : 325 ] * 11'b11111101001 + 
						X [ 348 : 337 ] * 11'b11111010011 + X [ 360 : 349 ] * 10'b1111110101 + 
						{X [ 372 : 361 ], 10'b0000000000} + X [ 384 : 373 ] * 11'b10111101111 + 
						X [ 396 : 385 ] * 12'b110111010011 + X [ 408 : 397 ] * 11'b10011110010 + 
						{X [ 420 : 409 ], 8'b00000000} + X [ 432 : 421 ] * 12'b110101011010 + 
						X [ 444 : 433 ] * 12'b111101010011 + X [ 456 : 445 ] * 12'b100100100110 + 
						{X [ 468 : 457 ], 6'b000000} + X [ 480 : 469 ] * 12'b101101000000 + 
						X [ 492 : 481 ] * 12'b111110110011 + X [ 500 : 493 ] * 12'b101000110011 ;

assign R_temp_2 = R_temp_1 [ 12 : 1 ]  + R_temp_1 [ 24 : 13 ] * 6'b101101 + 
						R_temp_1 [ 28 : 25 ] * 11'b11111101001 ;

assign R_temp_3 = R_temp_2 [ 12 : 1 ]  + R_temp_2 [18 : 13 ] * 6'b101101 ;

assign R_temp_4 = R_temp_3 [ 12 : 1 ]  + R_temp_3 [ 13 ] * 6'b101101 ;

always @(R_temp_4)
begin
  if (R_temp_4 >= 12'b111111010011)
    R_temp <= R_temp_4 - 12'b111111010011;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
