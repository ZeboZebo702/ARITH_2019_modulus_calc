module x_500_mod_461(
    input [500:1] X,
    output [9:1] R
    );

wire [23:1] R_temp_1;
wire [15:1] R_temp_2;
wire [12:1] R_temp_3;
wire [10:1] R_temp_4;
reg [9:1]  R_temp;

assign R_temp_1 = X [ 9 : 1 ]  + X [ 18 : 10 ] * 6'b110011 + X [ 27 : 19 ] * 9'b100101000 + X [ 36 : 28 ] * 9'b101011000 + X [ 45 : 37 ] * 5'b11010 + X [ 54 : 46 ] * 9'b110010100 + X [ 63 : 55 ] * 9'b101000000 + X [ 72 : 64 ] * 8'b10111001 + X [ 81 : 73 ] * 8'b11010111 + X [ 90 : 82 ] * 9'b101101010 + X [ 99 : 91 ] * 5'b10110 + X [ 108 : 100 ] * 8'b11001000 + X [ 117 : 109 ] * 6'b111010 + X [ 126 : 118 ] * 8'b11000000 + X [ 135 : 127 ] * 7'b1101111 + X [ 144 : 136 ] * 8'b10000001 + X [ 153 : 145 ] * 7'b1111101 + X [ 162 : 154 ] * 9'b101111110 + X [ 171 : 163 ] * 7'b1111000 + X [ 180 : 172 ] * 7'b1111111 + X [ 189 : 181 ] * 5'b10111 + X [ 198 : 190 ] * 8'b11111011 + X [ 207 : 199 ] * 9'b101100010 + X [ 216 : 208 ] * 7'b1001011 + X [ 225 : 217 ] * 8'b10001001 + X [ 234 : 226 ] * 7'b1001000 + X [ 243 : 235 ] * 9'b110111101 + X [ 252 : 244 ] * 7'b1101010 + X [ 261 : 253 ] * 9'b101001111 + X [ 270 : 262 ] * 5'b11100 + X [ 279 : 271 ] * 6'b101101 + X [ 288 : 280 ] * 9'b111000011 + X [ 297 : 289 ] * 9'b110011100 + X [ 306 : 298 ] * 9'b100001011 + X [ 315 : 307 ] * 8'b11111000 + X [ 324 : 316 ] * 8'b11001001 + X [ 333 : 325 ] * 7'b1101101 + X [ 342 : 334 ] * 5'b11011 + X [ 351 : 343 ] * 9'b111000111 + X [ 360 : 352 ] * 8'b10011011 + X [ 369 : 361 ] * 7'b1000100 + X [ 378 : 370 ] * 8'b11110001 + X [ 387 : 379 ] * 9'b100110001 + X [ 396 : 388 ] * 9'b101010110 + X [ 405 : 397 ] * 9'b110000001 + X [ 414 : 406 ] * 9'b100010001 + X [ 423 : 415 ] * 7'b1011101 + X [ 432 : 424 ] * 8'b10000101 + X [ 441 : 433 ] * 9'b101001001 + X [ 450 : 442 ] * 8'b10110111 + X [ 459 : 451 ] * 7'b1110001 + X [ 468 : 460 ] * 8'b11100111 + X [ 477 : 469 ] * 9'b100000000 + X [ 486 : 478 ] * 8'b10010100 + X [ 495 : 487 ] * 8'b10101100 + X [ 500 : 496 ] * 4'b1101 ;

assign R_temp_2 = R_temp_1 [ 9 : 1 ]  + R_temp_1 [ 18 : 10 ] * 6'b110011 + R_temp_1 [ 23 : 19 ] * 9'b100101000 ;

assign R_temp_3 = R_temp_2 [ 9 : 1 ]  + R_temp_2 [ 15 : 10 ] * 6'b110011 ;

assign R_temp_4 = R_temp_3 [ 9 : 1 ]  + R_temp_3 [ 12 :10 ] * 6'b110011 ;


always @(R_temp_4)
begin
  if (R_temp_4 >= 9'b111001101)
    R_temp <= R_temp_4 - 9'b111001101;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
