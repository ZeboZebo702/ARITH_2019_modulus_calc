module x_400_mod_107	(
    input [400:1] X,
    output [7:1] R
    );

wire [19:1] R_temp_1;
wire [12:1] R_temp_2;
wire [10:1] R_temp_3;
wire [8:1] R_temp_4;
reg [7:1]  R_temp;

assign R_temp_1 = X [ 7 : 1 ]  + X [ 14 : 8 ] * 5'b10101 + X [ 21 : 15 ] * 4'b1101 + X [ 28 : 22 ] * 6'b111011 + X [ 35 : 29 ] * 6'b111110 + 
		  X [ 42 : 36 ] * 5'b10010 + X [ 49 : 43 ] * 6'b111001 + X [ 56 : 50 ] * 5'b10100 + X [ 63 : 57 ] * 7'b1100011 + 
		  X [ 70 : 64 ] * 6'b101110 + X [ 77 : 71 ] * 2'b11 + X [ 84 : 78 ] * 6'b111111 + X [ 91 : 85 ] * 6'b100111 + 
		  X [ 98 : 92 ] * 7'b1000110 + X [ 105 : 99 ] * 7'b1001111 + X [ 112 : 106 ] * 6'b110110 + 
		  X [ 119 : 113 ] * 7'b1000000 + X [ 126 : 120 ] * 6'b111100 + X [ 133 : 127 ] * 7'b1010011 + X [ 140 : 134 ] * 5'b11111 + 
		  X [ 147 : 141 ] * 4'b1001 + X [ 154 : 148 ] * 7'b1010010 + X [ 161 : 155 ] * 4'b1010 + X [ 168 : 162 ] * 7'b1100111 + 
		  X [ 175 : 169 ] * 5'b10111 + X [ 182 : 176 ] * 6'b110111 + X [ 189 : 183 ] * 7'b1010101 + X [ 196 : 190 ] * 7'b1001001 + 
		  X [ 203 : 197 ] * 6'b100011 + X [ 210 : 204 ] * 7'b1011101 + X [ 217 : 211 ] * 5'b11011 + X [ 224 : 218 ] * 6'b100000 + 
		  X [ 231 : 225 ] * 5'b11110 + X [ 238 : 232 ] * 7'b1011111 + X [ 245 : 239 ] * 7'b1000101 + X [ 252 : 246 ] * 6'b111010 + 
		  X [ 259 : 253 ] * 6'b101001 + X [ 266 : 260 ] * 3'b101 + X [ 273 : 267 ] * 7'b1101001 + X [ 280 : 274 ] * 7'b1000001 + 
		  X [ 287 : 281 ] * 7'b1010001 + X [ 294 : 288 ] * 7'b1100000 + X [ 301 : 295 ] * 7'b1011010 + X [ 308 : 302 ] * 7'b1000111 + 
		  X [ 315 : 309 ] * 7'b1100100 + X [ 322 : 316 ] * 7'b1000011 + X [ 329 : 323 ] * 5'b10000 + X [ 336 : 330 ] * 4'b1111 + 
		  X [ 343 : 337 ] * 7'b1100101 + X [ 350 : 344 ] * 7'b1011000 + X [ 357 : 351 ] * 5'b11101 + X [ 364 : 358 ] * 7'b1001010 + 
		  X [ 371 : 365 ] * 6'b111000 + X [ 378 : 372 ] * 7'b1101010 + X [ 385 : 379 ] * 7'b1010110 + X [ 392 : 386 ] * 7'b1011110 + 
		  X [ 399 : 393 ] * 6'b110000 + X [ 400 ] * 6'b101101;

assign R_temp_2 = R_temp_1 [ 7 : 1 ]  + R_temp_1 [ 14 : 8 ] * 5'b10101 + R_temp_1 [ 19 : 15 ] * 4'b1101 ;

assign R_temp_3 = R_temp_2 [ 7 : 1 ]  + R_temp_2 [ 12 : 8 ] * 5'b10101 ;

assign R_temp_4 = R_temp_3 [ 7 : 1 ]  + R_temp_3 [ 10 : 8 ] * 5'b10101;

always @(R_temp_4)
begin
  if (R_temp_4 >= 7'b1101011)
    R_temp <= R_temp_4 - 7'b1101011;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
