module x_200_mod_107	(
    input [200:1] X,
    output [7:1] R
    );

wire [18:1] R_temp_1;
wire [12:1] R_temp_2;
wire [10:1] R_temp_3;
wire [8:1] R_temp_4;
reg [7:1]  R_temp;

assign R_temp_1 = X [ 7 : 1 ]  + X [ 14 : 8 ] * 5'b10101 + X [ 21 : 15 ] * 4'b1101 + X [ 28 : 22 ] * 6'b111011 + X [ 35 : 29 ] * 6'b111110 + 
		  X [ 42 : 36 ] * 5'b10010 + X [ 49 : 43 ] * 6'b111001 + X [ 56 : 50 ] * 5'b10100 + X [ 63 : 57 ] * 7'b1100011 + 
		  X [ 70 : 64 ] * 6'b101110 + X [ 77 : 71 ] * 2'b11 + X [ 84 : 78 ] * 6'b111111 + X [ 91 : 85 ] * 6'b100111 + 
		  X [ 98 : 92 ] * 7'b1000110 + X [ 105 : 99 ] * 7'b1001111 + X [ 112 : 106 ] * 6'b110110 + 
		  X [ 119 : 113 ] * 7'b1000000 + X [ 126 : 120 ] * 6'b111100 + X [ 133 : 127 ] * 7'b1010011 + X [ 140 : 134 ] * 5'b11111 + 
		  X [ 147 : 141 ] * 4'b1001 + X [ 154 : 148 ] * 7'b1010010 + X [ 161 : 155 ] * 4'b1010 + X [ 168 : 162 ] * 7'b1100111 + 
		  X [ 175 : 169 ] * 5'b10111 + X [ 182 : 176 ] * 6'b110111 + X [ 189 : 183 ] * 7'b1010101 + X [ 196 : 190 ] * 7'b1001001 + 
		  X [ 200 : 197 ] * 6'b100011 ;

assign R_temp_2 = R_temp_1 [ 7 : 1 ]  + R_temp_1 [ 14 : 8 ] * 5'b10101 + R_temp_1 [ 18 : 15 ] * 4'b1101 ;

assign R_temp_3 = R_temp_2 [ 7 : 1 ]  + R_temp_2 [ 12 : 8 ] * 5'b10101 ;

assign R_temp_4 = R_temp_3 [ 7 : 1 ]  + R_temp_3 [ 10 : 8 ] * 5'b10101;

always @(R_temp_4)
begin
  if (R_temp_4 >= 7'b1101011)
    R_temp <= R_temp_4 - 7'b1101011;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
