module x_300_mod_47(
    input [300:1] X,
    output [6:1] R
    );

wire [16:1] R_temp_1;
wire [11:1] R_temp_2;
wire [9:1] R_temp_3;
wire [8:1] R_temp_4;
wire [7:1] R_temp_5;
reg [6:1]  R_temp;

assign R_temp_1 = X [ 6 : 1 ]  + X [ 12 : 7 ] * 5'b10001 + X [ 18 : 13 ] * 3'b111 + X [ 24 : 19 ] * 5'b11001 + X [ 30 : 25 ] * 2'b10 + X [ 36 : 31 ] * 6'b100010 + X [ 42 : 37 ] * 4'b1110 + X [ 48 : 43 ] * 2'b11 + X [ 54 : 49 ] * 3'b100 + X [ 60 : 55 ] * 5'b10101 + X [ 66 : 61 ] * 5'b11100 + X [ 72 : 67 ] * 3'b110 + X [ 78 : 73 ] * 4'b1000 + X [ 84 : 79 ] * 6'b101010 + X [ 90 : 85 ] * 4'b1001 + X [ 96 : 91 ] * 4'b1100 + X [ 102 : 97 ] * 5'b10000 + X [ 108 : 103 ] * 6'b100101 + X [ 114 : 109 ] * 5'b10010 + X [ 120 : 115 ] * 5'b11000 + X [ 126 : 121 ] * 6'b100000 + X [ 132 : 127 ] * 5'b11011 + X [ 138 : 133 ] * 6'b100100 + X [ 144 : 139 ]  + X [ 150 : 145 ] * 5'b10001 + X [ 156 : 151 ] * 3'b111 + X [ 162 : 157 ] * 5'b11001 + X [ 168 : 163 ] * 2'b10 + X [ 174 : 169 ] * 6'b100010 + X [ 180 : 175 ] * 4'b1110 + X [ 186 : 181 ] * 2'b11 + X [ 192 : 187 ] * 3'b100 + X [ 198 : 193 ] * 5'b10101 + X [ 204 : 199 ] * 5'b11100 + X [ 210 : 205 ] * 3'b110 + X [ 216 : 211 ] * 4'b1000 + X [ 222 : 217 ] * 6'b101010 + X [ 228 : 223 ] * 4'b1001 + X [ 234 : 229 ] * 4'b1100 + X [ 240 : 235 ] * 5'b10000 + X [ 246 : 241 ] * 6'b100101 + X [ 252 : 247 ] * 5'b10010 + X [ 258 : 253 ] * 5'b11000 + X [ 264 : 259 ] * 6'b100000 + X [ 270 : 265 ] * 5'b11011 + X [ 276 : 271 ] * 6'b100100 + X [ 282 : 277 ]  + X [ 288 : 283 ] * 5'b10001 + X [ 294 : 289 ] * 3'b111 + X [ 300 : 295 ] * 5'b11001 ;

assign R_temp_2 = R_temp_1 [6 : 1]  + R_temp_1 [ 12 : 7 ] * 5'b10001 + R_temp_1 [ 16 : 13 ] * 3'b111 ;

assign R_temp_3 = R_temp_2 [6 : 1]  + R_temp_2 [ 11 : 7 ] * 5'b10001;

assign R_temp_4 = R_temp_3 [6 : 1]  + R_temp_3 [ 9 : 7 ] * 5'b10001;

assign R_temp_5 = R_temp_4 [6 : 1]  + R_temp_4 [ 8 : 7 ] * 5'b10001;

always @(R_temp_5)
begin
  if (R_temp_5 >= 6'b101111)
    R_temp <= R_temp_5 - 6'b101111;
  else
    R_temp <= R_temp_5;
end

assign R = R_temp;

endmodule
