module x_300_mod_4051(
    input [300:1] X,
    output [12:1] R
    );

wire [28:1] R_temp_1;
wire [18:1] R_temp_2;
wire [13:1] R_temp_3;
wire [13:1] R_temp_4;
reg [12:1]  R_temp;

assign R_temp_1 = X [ 12 : 1 ]  + X [ 24 : 13 ] * 6'b101101 + X [ 36 : 25 ] * 11'b11111101001 + 
						X [ 48 : 37 ] * 11'b11111010011 + X [ 60 : 49 ] * 10'b1111110101 + 
						{X [ 72 : 61 ], 10'b0000000000} + X [ 84 : 73 ] * 11'b10111101111 + 
						X [ 96 : 85 ] * 12'b110111010011 + X [ 108 : 97 ] * 11'b10011110010 + 
						{X [ 120 : 109 ], 8'b00000000} + X [ 132 : 121 ] * 12'b110101011010 + 
						X [ 144 : 133 ] * 12'b111101010011 + X [ 156 : 145 ] * 12'b100100100110 + 
						{X [ 168 : 157 ], 6'b000000} + X [ 180 : 169 ] * 12'b101101000000 + 
						X [ 192 : 181 ] * 12'b111110110011 + X [ 204 : 193 ] * 12'b101000110011 + 
						{X [ 216 : 205 ], 4'b0000} + X [ 228 : 217 ] * 10'b1011010000 + 
						X [ 240 : 229 ] * 12'b111111001011 + X [ 252 : 241 ] * 12'b111001101011 + 
						{X [ 264 : 253 ], 2'b00} + X [ 276 : 265 ] * 8'b10110100 + 
						X [ 288 : 277 ] * 12'b111111010001 + X [ 300 : 289 ] * 12'b111101111001 ;

assign R_temp_2 = R_temp_1 [ 12 : 1 ]  + R_temp_1 [ 24 : 13 ] * 6'b101101 + 
						R_temp_1 [ 28 : 25 ] * 11'b11111101001 ;

assign R_temp_3 = R_temp_2 [ 12 : 1 ]  + R_temp_2 [18 : 13 ] * 6'b101101 ;

assign R_temp_4 = R_temp_3 [ 12 : 1 ]  + R_temp_3 [ 13 ] * 6'b101101 ;

always @(R_temp_4)
begin
  if (R_temp_4 >= 12'b111111010011)
    R_temp <= R_temp_4 - 12'b111111010011;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
