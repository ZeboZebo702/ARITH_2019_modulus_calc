module x_500_mod_53(
    input [500:1] X,
    output [6:1] R
    );

wire [18:1] R_temp_1;
wire [11:1] R_temp_2;
wire [8:1] R_temp_3;
wire [7:1] R_temp_4;
reg [6:1]  R_temp;

assign R_temp_1 = X [ 6 : 1 ]  + X [ 12 : 7 ] * 4'b1011 + X [ 18 : 13 ] * 4'b1111 + X [ 24 : 19 ] * 3'b110 + 
X [ 30 : 25 ] * 4'b1101 + X [ 36 : 31 ] * 6'b100101 + X [ 42 : 37 ] * 6'b100100 + X [ 48 : 43 ] * 5'b11001 + 
X [ 54 : 49 ] * 4'b1010 + {X [ 60 : 55 ], 2'b00} + X [ 66 : 61 ] * 6'b101100 + X [ 72 : 67 ] * 3'b111 + 
X [ 78 : 73 ] * 5'b11000 + X [ 84 : 79 ] * 6'b110100 + X [ 90 : 85 ] * 6'b101010 + X [ 96 : 91 ] * 6'b100110 + 
X [ 102 : 97 ] * 6'b101111 + X [ 108 : 103 ] * 6'b101000 + X [ 114 : 109 ] * 5'b10000 + 
X [ 120 : 115 ] * 5'b10001 + X [ 126 : 121 ] * 5'b11100 + X [ 132 : 127 ] * 6'b101011 + 
X [ 138 : 133 ] * 6'b110001 + X [ 144 : 139 ] * 4'b1001 + X [ 150 : 145 ] * 6'b101110 + 
X [ 156 : 151 ] * 5'b11101 + X [ 162 : 157 ]  + X [ 168 : 163 ] * 4'b1011 + X [ 174 : 169 ] * 4'b1111 + 
X [ 180 : 175 ] * 3'b110 + X [ 186 : 181 ] * 4'b1101 + X [ 192 : 187 ] * 6'b100101 + 
X [ 198 : 193 ] * 6'b100100 + X [ 204 : 199 ] * 5'b11001 + X [ 210 : 205 ] * 4'b1010 + 
{X [ 216 : 211 ], 2'b00} + X [ 222 : 217 ] * 6'b101100 + X [ 228 : 223 ] * 3'b111 + 
X [ 234 : 229 ] * 5'b11000 + X [ 240 : 235 ] * 6'b110100 + X [ 246 : 241 ] * 6'b101010 + 
X [ 252 : 247 ] * 6'b100110 + X [ 258 : 253 ] * 6'b101111 + X [ 264 : 259 ] * 6'b101000 + 
{X [ 270 : 265 ], 4'b0000} + X [ 276 : 271 ] * 5'b10001 + X [ 282 : 277 ] * 5'b11100 + 
X [ 288 : 283 ] * 6'b101011 + X [ 294 : 289 ] * 6'b110001 + X [ 300 : 295 ] * 4'b1001 + 
X [ 306 : 301 ] * 6'b101110 + X [ 312 : 307 ] * 5'b11101 + X [ 318 : 313 ]  + X [ 324 : 319 ] * 4'b1011 + 
X [ 330 : 325 ] * 4'b1111 + X [ 336 : 331 ] * 3'b110 + X [ 342 : 337 ] * 4'b1101 + 
X [ 348 : 343 ] * 6'b100101 + X [ 354 : 349 ] * 6'b100100 + X [ 360 : 355 ] * 5'b11001 + 
X [ 366 : 361 ] * 4'b1010 + {X [ 372 : 367 ], 2'b00} + X [ 378 : 373 ] * 6'b101100 + 
X [ 384 : 379 ] * 3'b111 + X [ 390 : 385 ] * 5'b11000 + X [ 396 : 391 ] * 6'b110100 + 
X [ 402 : 397 ] * 6'b101010 + X [ 408 : 403 ] * 6'b100110 + X [ 414 : 409 ] * 6'b101111 + 
X [ 420 : 415 ] * 6'b101000 + {X [ 426 : 421 ], 4'b0000} + X [ 432 : 427 ] * 5'b10001 + 
X [ 438 : 433 ] * 5'b11100 + X [ 444 : 439 ] * 6'b101011 + X [ 450 : 445 ] * 6'b110001 + 
X [ 456 : 451 ] * 4'b1001 + X [ 462 : 457 ] * 6'b101110 + X [ 468 : 463 ] * 5'b11101 + 
X [ 474 : 469 ]  + X [ 480 : 475 ] * 4'b1011 + X [ 486 : 481 ] * 4'b1111 + X [ 492 : 487 ] * 3'b110 + 
X [ 498 : 493 ] * 4'b1101 + X [ 500 : 499 ] * 6'b100101 ;

assign R_temp_2 = R_temp_1 [ 6 : 1 ]  + R_temp_1 [ 12 : 7 ] * 4'b1011 + R_temp_1 [ 18 : 13 ] * 4'b1111 ;

assign R_temp_3 = R_temp_2 [ 6 : 1 ]  + R_temp_2 [ 11 : 7 ] * 4'b1011 ;

assign R_temp_4 = R_temp_3 [ 6 : 1 ]  + R_temp_3 [ 8 : 7 ] * 4'b1011 ;

always @(R_temp_4)
begin
  if (R_temp_4 >= 6'b110101)
    R_temp <= R_temp_4 - 6'b110101;
  else
    R_temp <= R_temp_4;
end

assign R = R_temp;

endmodule
