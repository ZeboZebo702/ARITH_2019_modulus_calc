module x_500_mod_503(
    input [500:1] X,
    output [9:1] R
    );

wire [23:1] R_temp_1;
wire [13:1] R_temp_2;
wire [10:1] R_temp_3;
reg [9:1]  R_temp;

assign R_temp_1 =X [ 9 : 1 ]  + X [ 18 : 10 ] * 4'b1001 + X [ 27 : 19 ] * 7'b1010001 + 
X [ 36 : 28 ] * 8'b11100010 + X [ 45 : 37 ] * 5'b10110 + X [ 54 : 46 ] * 8'b11000110 + 
X [ 63 : 55 ] * 9'b100010001 + X [ 72 : 64 ] * 9'b110111101 + X [ 81 : 73 ] * 9'b111100100 + 
X [ 90 : 82 ] * 9'b101001100 + X [ 99 : 91 ] * 9'b111011001 + X [ 108 : 100 ] * 8'b11101001 + 
X [ 117 : 109 ] * 7'b1010101 + X [ 126 : 118 ] * 9'b100000110 + X [ 135 : 127 ] * 9'b101011010 + 
X [ 144 : 136 ] * 7'b1100000 + X [ 153 : 145 ] * 9'b101101001 + X [ 162 : 154 ] * 8'b11100111 + 
X [ 171 : 163 ] * 7'b1000011 + X [ 180 : 172 ] * 7'b1100100 + X [ 189 : 181 ] * 9'b110001101 + 
X [ 198 : 190 ] * 6'b110100 + X [ 207 : 199 ] * 9'b111010100 + X [ 216 : 208 ] * 8'b10111100 + 
X [ 225 : 217 ] * 8'b10110111 + X [ 234 : 226 ] * 8'b10001010 + X [ 243 : 235 ] * 8'b11101100 + 
X [ 252 : 244 ] * 7'b1110000 + X [ 261 : 253 ] * 2'b10 + X [ 270 : 262 ] * 5'b10010 + 
X [ 279 : 271 ] * 8'b10100010 + X [ 288 : 280 ] * 9'b111000100 + X [ 297 : 289 ] * 6'b101100 + 
X [ 306 : 298 ] * 9'b110001100 + X [ 315 : 307 ] * 6'b101011 + X [ 324 : 316 ] * 9'b110000011 + 
X [ 333 : 325 ] * 9'b111010001 + X [ 342 : 334 ] * 8'b10100001 + X [ 351 : 343 ] * 9'b110111011 + 
X [ 360 : 352 ] * 9'b111010010 + X [ 369 : 361 ] * 8'b10101010 + X [ 378 : 370 ] * 5'b10101 + 
X [ 387 : 379 ] * 8'b10111101 + X [ 396 : 388 ] * 8'b11000000 + X [ 405 : 397 ] * 8'b11011011 + 
X [ 414 : 406 ] * 9'b111001110 + X [ 423 : 415 ] * 8'b10000110 + X [ 432 : 424 ] * 8'b11001000 + 
X [ 441 : 433 ] * 9'b100100011 + X [ 450 : 442 ] * 7'b1101000 + X [ 459 : 451 ] * 9'b110110001 + 
X [ 468 : 460 ] * 9'b101111000 + X [ 477 : 469 ] * 9'b101101110 + X [ 486 : 478 ] * 9'b100010100 + 
X [ 495 : 487 ] * 9'b111011000 + X [ 500 : 496 ] * 8'b11100000 ;

assign R_temp_2 = R_temp_1 [ 9 : 1 ]  + R_temp_1 [ 18 : 10 ] * 4'b1001 + R_temp_1 [ 23 : 19 ] * 7'b1010001 ;

assign R_temp_3 = R_temp_2 [ 9 : 1 ]  + R_temp_2 [ 13 : 10 ] * 4'b1001 ;

always @(R_temp_3)
begin
  if (R_temp_3 >= 9'b111110111)
    R_temp <= R_temp_3 - 9'b111110111;
  else
    R_temp <= R_temp_3;
end

assign R = R_temp;

endmodule
